// Copyright (c) 2024 Andrew Parker

package env_pkg;

   import uvm_pkg::*;
`include "uvm_macros.svh"

   // Register bus agent
`include "reg_bus_item.svh"
`include "reg_bus_monitor.svh"
`include "reg_bus_driver.svh"
`include "reg_bus_agent.svh"
`include "reg_bus_seq_lib.svh"

   // Register model
`include "reg_model.svh"

   // Env
`include "env.svh"

endpackage: env_pkg
