// Copyright (c) 2024 Andrew Parker

package env_pkg;

   import uvm_pkg::*;
`include "uvm_macros.svh"

   // Reg agent
`include "reg_item.svh"
`include "reg_monitor.svh"
`include "reg_driver.svh"
`include "reg_agent.svh"
`include "reg_seq_lib.svh"

   // Env
`include "env.svh"

endpackage: env_pkg
