// Copyright (c) 2024 Andrew Parker

package test_pkg;

   import uvm_pkg::*;
`include "uvm_macros.svh"

endpackage: test_pkg
